`timescale 1ns / 1ps

interface dff_if();

bit clk;
bit rst;
logic din;
logic dout;

endinterface
